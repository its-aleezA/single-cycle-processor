//OR gate module
module OR(a, b, c);
    input a, b;
    output c;
    
    assign c = a | b;
endmodule
